BZh91AY&SYq�1  �_�Px���g߰?���@v��mWs�(��jz��LOH�h�S�44 @��	"j�(��hOS��A�!����i�z�A�       SQ��@�I���j����   �F�qHE� í͌(�e���� �Q�i� ކ�x��tYe�������T@��Kc�<DW QQ�I�ET�5�++'C*�V�յ���"^.ANx����⦌�MC�VG
��ʩ1��6ʻV����86�0��T�טx���lhI��"3VhkC���A;�Q~I��Q���b;"�
��m��ǯ���2����H���w��&�=�]��#�̢��֛�J��/�,����eɬ�����K�ea�EG�`GbT��ppYHi�vsF�Օ����Dh�Z�f����|�^L�Y�D�U:X�l
�M!|$�
LH�!��ad���\t�i"_$��]Ár�*^��S&P�.&3�I�i`@]ah#/�AAy�C�5 �ptH
GT
K䴪aAF��K��&Y��X�ldG�J�af�E���Ӷ�aT�)`�����8"0�P��̸�m�XѤ��r�J���'�^�c�͔�#v���7/ZE*�1⡇�C�S�d��w�"_���w$S�	�S